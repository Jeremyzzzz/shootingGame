/***************************************************
module	:seg7_decoder
input	:��λ��Ҫ�����BCD��
output	:�߶�����ܵĶ������
function:��DE2��������ʵ����4λ���������

***************************************************/
module seg7_decoder(
	dat1_i,
	dat2_i,
	dat3_i,
	dat4_i,
	seg1_o,
	seg2_o,
	seg3_o,
	seg4_o
	); 

	input	[3:0]	dat1_i;				//��1λҪ��ʾ������
	input	[3:0]	dat2_i;				//��2λҪ��ʾ������
	input	[3:0]	dat3_i;				//��3λҪ��ʾ������
	input	[3:0]	dat4_i;				//��4λҪ��ʾ������
	
	output	[6:0]	seg1_o;				//��1λ�����������		
	output	[6:0]	seg2_o;				//��2λ�����������
	output	[6:0]	seg3_o;				//��3λ�����������
	output	[6:0]	seg4_o;				//��4λ�����������
	
	//����Ĵ�������								
	reg		[6:0]	seg1_o;				
	reg		[6:0]	seg2_o;				
	reg		[6:0]	seg3_o;				
	reg		[6:0]	seg4_o;
	
	always @(*)begin
		case(dat1_i)				//��1λ�����߶�����	
	//---------------------------------����-----------------------------------//	
			4'h0:seg1_o=7'b1000000;	//��ʾ0
			4'h1:seg1_o=7'b1111001;	//��ʾ1
			4'h2:seg1_o=7'b0100100;	//��ʾ2
			4'h3:seg1_o=7'b0110000;	//��ʾ3
			4'h4:seg1_o=7'b0011001;	//��ʾ4
			4'h5:seg1_o=7'b0010010;	//��ʾ5
			4'h6:seg1_o=7'b0000010;	//��ʾ6
			4'h7:seg1_o=7'b1111000;	//��ʾ7
			4'h8:seg1_o=7'b0000000;	//��ʾ8
			4'h9:seg1_o=7'b0011000;	//��ʾ9		
			default:seg1_o=7'b1111111;//����ʾ
		endcase
	end

	always @(*)begin
		case(dat2_i)				//��2λ�����߶�����	
	//---------------------------------����-----------------------------------//	
			4'h0:seg2_o=7'b1000000;	//��ʾ0
			4'h1:seg2_o=7'b1111001;	//��ʾ1
			4'h2:seg2_o=7'b0100100;	//��ʾ2
			4'h3:seg2_o=7'b0110000;	//��ʾ3
			4'h4:seg2_o=7'b0011001;	//��ʾ4
			4'h5:seg2_o=7'b0010010;	//��ʾ5
			4'h6:seg2_o=7'b0000010;	//��ʾ6
			4'h7:seg2_o=7'b1111000;	//��ʾ7
			4'h8:seg2_o=7'b0000000;	//��ʾ8
			4'h9:seg2_o=7'b0011000;	//��ʾ9
			default:seg2_o=7'b1111111;//����ʾ
		endcase
	end

	always @(*)begin
		case(dat3_i)				//��3λ�����߶�����	
	//---------------------------------����-----------------------------------//	
			4'h0:seg3_o=7'b1000000;	//��ʾ0
			4'h1:seg3_o=7'b1111001;	//��ʾ1
			4'h2:seg3_o=7'b0100100;	//��ʾ2
			4'h3:seg3_o=7'b0110000;	//��ʾ3
			4'h4:seg3_o=7'b0011001;	//��ʾ4
			4'h5:seg3_o=7'b0010010;	//��ʾ5
			4'h6:seg3_o=7'b0000010;	//��ʾ6
			4'h7:seg3_o=7'b1111000;	//��ʾ7
			4'h8:seg3_o=7'b0000000;	//��ʾ8
			4'h9:seg3_o=7'b0011000;	//��ʾ9
			default:seg3_o=7'b1111111;//����ʾ
		endcase
	end

	always @(*)begin
		case(dat4_i)				//��4λ�����߶�����	
	//---------------------------------����-----------------------------------//	
			4'h0:seg4_o=7'b1000000;	//��ʾ0
			4'h1:seg4_o=7'b1111001;	//��ʾ1
			4'h2:seg4_o=7'b0100100;	//��ʾ2
			4'h3:seg4_o=7'b0110000;	//��ʾ3
			4'h4:seg4_o=7'b0011001;	//��ʾ4
			4'h5:seg4_o=7'b0010010;	//��ʾ5
			4'h6:seg4_o=7'b0000010;	//��ʾ6
			4'h7:seg4_o=7'b1111000;	//��ʾ7
			4'h8:seg4_o=7'b0000000;	//��ʾ8
			4'h9:seg4_o=7'b0011000;	//��ʾ9		
			default:seg4_o=7'b1111111;//����ʾ
		endcase
	end
	
endmodule
